//
// Verilog Module encoder_decoder_lib.ECC_ENC_DEC
//
// Created:
//          by - yuvalsaa.UNKNOWN (L330W530)
//          at - 15:59:09 11/10/2021
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module ECC_ENC_DEC ;


// ### Please start your Verilog code here ### 

endmodule
