//
// Verilog Module encoder_decoder_lib.dec_is_column
//
// Created:
//          by - yuvalsaa.UNKNOWN (L330W530)
//          at - 17:41:52 11/10/2021
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module dec_is_column ;


// ### Please start your Verilog code here ### 

endmodule
