//
// Verilog Module encoder_decoder_lib.enc_parity_16bit
//
// Created:
//          by - yuvalsaa.UNKNOWN (L330W530)
//          at - 17:33:17 11/10/2021
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module enc_parity_16bit ;


// ### Please start your Verilog code here ### 

endmodule
