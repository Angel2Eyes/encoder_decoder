//
// Verilog Module encoder_decoder_lib.verification_checker
//
// Created:
//          by - yuvalsaa.UNKNOWN (L330W527)
//          at - 15:00:13 12/19/2021
//
// using Mentor Graphics HDL Designer(TM) 2016.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module verification_checker ;


// ### Please start your Verilog code here ### 

endmodule
